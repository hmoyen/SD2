module datapath (clock, a, b, sinal, state, res);


    input wire [3:0] state;
    reg [4:0] num1, num2;
    reg [15:0] num3, num4;
    reg [15:0] some, someXYShift;
    reg [8:0] someXY;
    reg [9:0] subDEXY;
    reg [13:0] subShift;
    reg [9:0] produtoDE;
    reg [7:0] X, Y;
    reg [8:0] A;
    reg [8:0] B;
    output reg [16:0] res;
    reg [4:0] E, D;
    reg [15:0] shiftY;
    reg[3:0] aH, bH, aL, bL;
    input [8:0] a;
    input [8:0] b;
    output reg [9:0] z;
    reg mag_a, mag_b, mag_res;
    input wire clock, start;
    input sinal;
    parameter IDLE = 4'b0000, MUL0 = 4'b0001, MUL1 = 4'b0010, MUL2 = 4'b0011,
    MUL3 = 4'b0100, MUL4 = 4'b0101, MUL5 = 4'b0110, MUL6 = 4'b0111, MUL7 = 4'b1000, MUL8 = 4'b1001, MUL9 = 4'b1010, DONE = 4'b1011;

    always@(posedge clock)
    begin

        case(state)

            IDLE:
            begin
                
                A <= ~(a - 1'b1);
                $display("%b",A);
                B <= ~(b - 1'b1);
                $display("%b",B);

                
                
                // $display("%b",a);
                

                res <=0;
                X <= 0;
                Y <= 0;
                E <= 0;
                D <= 0;

                someXY <= 0;
                someXYShift <= 0;
                subDEXY <= 0;
                subShift <=0;
                shiftY <= 0;
                produtoDE <=0;
                
            end

            MUL0:
                begin
                    aH = A[7:4];
                    aL = A[3:0];
                    bH = B[7:4];
                    bL = B[3:0];
                    num1 <= aL;
                    num2 <= bL;
                    num3 <= bH;
                    num4 <= bL;
                    mag_a = A[8:8];
                    mag_b = B[8:8];
                    if (mag_a == mag_b)
                        mag_res = 0;
                    else 
                        mag_res = 1;
                end


            MUL1:
                begin
            
                    $display("%b",A);
                    X <= z;
                    E <= some;
                    
                    num1 <= aH;
                    num2 <= bH;
                    num3 <= aH;
                    num4 <= aL;
                    
                    
                end
            MUL2:
                begin
                    $display("%b", A);
                    Y <= z; 
                    D <= some;
                    
                    
                end
            MUL3:
                begin
                    
                    num1 <= D;
                    num2 <= E;
                    num3 <=X;
                    num4 <= Y;
                
                    
                    
                
                end
            MUL4:
                begin
                    someXY <= some;
                    produtoDE <= z;
            
                    
                end
            
            MUL5:
                begin
                    num3 <= produtoDE;
                    num4 <= someXY;
                    shiftY <= Y<<8;
                   
                end
            
            MUL6:
                begin
                    subDEXY <= some;
                    
                    num3 <= X;
                    num4 <= shiftY;
                    
                end
                    
            
            MUL7:
                begin
                    subShift <= subDEXY<<4;
                    someXYShift <= some;
                    
        
                end
            
            MUL8:
                begin
                    
                    num3 <= someXYShift;
                    num4 <= subShift;
                  
                    
                end
            
            MUL9:
                begin
                    res <= ~(some + 1'b1);
                    res[16:16] <= mag_res;

                    
                end
            DONE:
                begin
                    
                    $display("%b",res);
                    $finish;
                end
                


            
  
        endcase
        end


    always @(num3,num4) begin

        
        if (sinal == 1'b0)
        begin

            some = num3 + num4;
            
           
            
        end
        else
        begin
            some = num3 - num4;
          
        end
        end
    

    always @(num1, num2) begin

        case ({num1, num2})
            10'b0000000000: z <= 10'b0000000000; // 0 * 0 = 0
            10'b0000000001: z <= 10'b0000000000; // 0 * 1 = 0
            10'b0000000010: z <= 10'b0000000000; // 0 * 2 = 0
            10'b0000000011: z <= 10'b0000000000; // 0 * 3 = 0
            10'b0000000100: z <= 10'b0000000000; // 0 * 4 = 0
            10'b0000000101: z <= 10'b0000000000; // 0 * 5 = 0
            10'b0000000110: z <= 10'b0000000000; // 0 * 6 = 0
            10'b0000000111: z <= 10'b0000000000; // 0 * 7 = 0
            10'b0000001000: z <= 10'b0000000000; // 0 * 8 = 0
            10'b0000001001: z <= 10'b0000000000; // 0 * 9 = 0
            10'b0000001010: z <= 10'b0000000000; // 0 * 10 = 0
            10'b0000001011: z <= 10'b0000000000; // 0 * 11 = 0
            10'b0000001100: z <= 10'b0000000000; // 0 * 12 = 0
            10'b0000001101: z <= 10'b0000000000; // 0 * 13 = 0
            10'b0000001110: z <= 10'b0000000000; // 0 * 14 = 0
            10'b0000001111: z <= 10'b0000000000; // 0 * 15 = 0
            10'b0000010000: z <= 10'b0000000000; // 0 * 16 = 0
            10'b0000010001: z <= 10'b0000000000; // 0 * 17 = 0
            10'b0000010010: z <= 10'b0000000000; // 0 * 18 = 0
            10'b0000010011: z <= 10'b0000000000; // 0 * 19 = 0
            10'b0000010100: z <= 10'b0000000000; // 0 * 20 = 0
            10'b0000010101: z <= 10'b0000000000; // 0 * 21 = 0
            10'b0000010110: z <= 10'b0000000000; // 0 * 22 = 0
            10'b0000010111: z <= 10'b0000000000; // 0 * 23 = 0
            10'b0000011000: z <= 10'b0000000000; // 0 * 24 = 0
            10'b0000011001: z <= 10'b0000000000; // 0 * 25 = 0
            10'b0000011010: z <= 10'b0000000000; // 0 * 26 = 0
            10'b0000011011: z <= 10'b0000000000; // 0 * 27 = 0
            10'b0000011100: z <= 10'b0000000000; // 0 * 28 = 0
            10'b0000011101: z <= 10'b0000000000; // 0 * 29 = 0
            10'b0000011110: z <= 10'b0000000000; // 0 * 30 = 0
            10'b0000011111: z <= 10'b0000000000; // 0 * 31 = 0
            10'b0000100000: z <= 10'b0000000000; // 1 * 0 = 0
            10'b0000100001: z <= 10'b0000000001; // 1 * 1 = 1
            10'b0000100010: z <= 10'b0000000010; // 1 * 2 = 2
            10'b0000100011: z <= 10'b0000000011; // 1 * 3 = 3
            10'b0000100100: z <= 10'b0000000100; // 1 * 4 = 4
            10'b0000100101: z <= 10'b0000000101; // 1 * 5 = 5
            10'b0000100110: z <= 10'b0000000110; // 1 * 6 = 6
            10'b0000100111: z <= 10'b0000000111; // 1 * 7 = 7
            10'b0000101000: z <= 10'b0000001000; // 1 * 8 = 8
            10'b0000101001: z <= 10'b0000001001; // 1 * 9 = 9
            10'b0000101010: z <= 10'b0000001010; // 1 * 10 = 10
            10'b0000101011: z <= 10'b0000001011; // 1 * 11 = 11
            10'b0000101100: z <= 10'b0000001100; // 1 * 12 = 12
            10'b0000101101: z <= 10'b0000001101; // 1 * 13 = 13
            10'b0000101110: z <= 10'b0000001110; // 1 * 14 = 14
            10'b0000101111: z <= 10'b0000001111; // 1 * 15 = 15
            10'b0000110000: z <= 10'b0000010000; // 1 * 16 = 16
            10'b0000110001: z <= 10'b0000010001; // 1 * 17 = 17
            10'b0000110010: z <= 10'b0000010010; // 1 * 18 = 18
            10'b0000110011: z <= 10'b0000010011; // 1 * 19 = 19
            10'b0000110100: z <= 10'b0000010100; // 1 * 20 = 20
            10'b0000110101: z <= 10'b0000010101; // 1 * 21 = 21
            10'b0000110110: z <= 10'b0000010110; // 1 * 22 = 22
            10'b0000110111: z <= 10'b0000010111; // 1 * 23 = 23
            10'b0000111000: z <= 10'b0000011000; // 1 * 24 = 24
            10'b0000111001: z <= 10'b0000011001; // 1 * 25 = 25
            10'b0000111010: z <= 10'b0000011010; // 1 * 26 = 26
            10'b0000111011: z <= 10'b0000011011; // 1 * 27 = 27
            10'b0000111100: z <= 10'b0000011100; // 1 * 28 = 28
            10'b0000111101: z <= 10'b0000011101; // 1 * 29 = 29
            10'b0000111110: z <= 10'b0000011110; // 1 * 30 = 30
            10'b0000111111: z <= 10'b0000011111; // 1 * 31 = 31
            10'b0001000000: z <= 10'b0000000000; // 2 * 0 = 0
            10'b0001000001: z <= 10'b0000000010; // 2 * 1 = 2
            10'b0001000010: z <= 10'b0000000100; // 2 * 2 = 4
            10'b0001000011: z <= 10'b0000000110; // 2 * 3 = 6
            10'b0001000100: z <= 10'b0000001000; // 2 * 4 = 8
            10'b0001000101: z <= 10'b0000001010; // 2 * 5 = 10
            10'b0001000110: z <= 10'b0000001100; // 2 * 6 = 12
            10'b0001000111: z <= 10'b0000001110; // 2 * 7 = 14
            10'b0001001000: z <= 10'b0000010000; // 2 * 8 = 16
            10'b0001001001: z <= 10'b0000010010; // 2 * 9 = 18
            10'b0001001010: z <= 10'b0000010100; // 2 * 10 = 20
            10'b0001001011: z <= 10'b0000010110; // 2 * 11 = 22
            10'b0001001100: z <= 10'b0000011000; // 2 * 12 = 24
            10'b0001001101: z <= 10'b0000011010; // 2 * 13 = 26
            10'b0001001110: z <= 10'b0000011100; // 2 * 14 = 28
            10'b0001001111: z <= 10'b0000011110; // 2 * 15 = 30
            10'b0001010000: z <= 10'b0000100000; // 2 * 16 = 32
            10'b0001010001: z <= 10'b0000100010; // 2 * 17 = 34
            10'b0001010010: z <= 10'b0000100100; // 2 * 18 = 36
            10'b0001010011: z <= 10'b0000100110; // 2 * 19 = 38
            10'b0001010100: z <= 10'b0000101000; // 2 * 20 = 40
            10'b0001010101: z <= 10'b0000101010; // 2 * 21 = 42
            10'b0001010110: z <= 10'b0000101100; // 2 * 22 = 44
            10'b0001010111: z <= 10'b0000101110; // 2 * 23 = 46
            10'b0001011000: z <= 10'b0000110000; // 2 * 24 = 48
            10'b0001011001: z <= 10'b0000110010; // 2 * 25 = 50
            10'b0001011010: z <= 10'b0000110100; // 2 * 26 = 52
            10'b0001011011: z <= 10'b0000110110; // 2 * 27 = 54
            10'b0001011100: z <= 10'b0000111000; // 2 * 28 = 56
            10'b0001011101: z <= 10'b0000111010; // 2 * 29 = 58
            10'b0001011110: z <= 10'b0000111100; // 2 * 30 = 60
            10'b0001011111: z <= 10'b0000111110; // 2 * 31 = 62
            10'b0001100000: z <= 10'b0000000000; // 3 * 0 = 0
            10'b0001100001: z <= 10'b0000000011; // 3 * 1 = 3
            10'b0001100010: z <= 10'b0000000110; // 3 * 2 = 6
            10'b0001100011: z <= 10'b0000001001; // 3 * 3 = 9
            10'b0001100100: z <= 10'b0000001100; // 3 * 4 = 12
            10'b0001100101: z <= 10'b0000001111; // 3 * 5 = 15
            10'b0001100110: z <= 10'b0000010010; // 3 * 6 = 18
            10'b0001100111: z <= 10'b0000010101; // 3 * 7 = 21
            10'b0001101000: z <= 10'b0000011000; // 3 * 8 = 24
            10'b0001101001: z <= 10'b0000011011; // 3 * 9 = 27
            10'b0001101010: z <= 10'b0000011110; // 3 * 10 = 30
            10'b0001101011: z <= 10'b0000100001; // 3 * 11 = 33
            10'b0001101100: z <= 10'b0000100100; // 3 * 12 = 36
            10'b0001101101: z <= 10'b0000100111; // 3 * 13 = 39
            10'b0001101110: z <= 10'b0000101010; // 3 * 14 = 42
            10'b0001101111: z <= 10'b0000101101; // 3 * 15 = 45
            10'b0001110000: z <= 10'b0000110000; // 3 * 16 = 48
            10'b0001110001: z <= 10'b0000110011; // 3 * 17 = 51
            10'b0001110010: z <= 10'b0000110110; // 3 * 18 = 54
            10'b0001110011: z <= 10'b0000111001; // 3 * 19 = 57
            10'b0001110100: z <= 10'b0000111100; // 3 * 20 = 60
            10'b0001110101: z <= 10'b0000111111; // 3 * 21 = 63
            10'b0001110110: z <= 10'b0001000010; // 3 * 22 = 66
            10'b0001110111: z <= 10'b0001000101; // 3 * 23 = 69
            10'b0001111000: z <= 10'b0001001000; // 3 * 24 = 72
            10'b0001111001: z <= 10'b0001001011; // 3 * 25 = 75
            10'b0001111010: z <= 10'b0001001110; // 3 * 26 = 78
            10'b0001111011: z <= 10'b0001010001; // 3 * 27 = 81
            10'b0001111100: z <= 10'b0001010100; // 3 * 28 = 84
            10'b0001111101: z <= 10'b0001010111; // 3 * 29 = 87
            10'b0001111110: z <= 10'b0001011010; // 3 * 30 = 90
            10'b0001111111: z <= 10'b0001011101; // 3 * 31 = 93
            10'b0010000000: z <= 10'b0000000000; // 4 * 0 = 0
            10'b0010000001: z <= 10'b0000000100; // 4 * 1 = 4
            10'b0010000010: z <= 10'b0000001000; // 4 * 2 = 8
            10'b0010000011: z <= 10'b0000001100; // 4 * 3 = 12
            10'b0010000100: z <= 10'b0000010000; // 4 * 4 = 16
            10'b0010000101: z <= 10'b0000010100; // 4 * 5 = 20
            10'b0010000110: z <= 10'b0000011000; // 4 * 6 = 24
            10'b0010000111: z <= 10'b0000011100; // 4 * 7 = 28
            10'b0010001000: z <= 10'b0000100000; // 4 * 8 = 32
            10'b0010001001: z <= 10'b0000100100; // 4 * 9 = 36
            10'b0010001010: z <= 10'b0000101000; // 4 * 10 = 40
            10'b0010001011: z <= 10'b0000101100; // 4 * 11 = 44
            10'b0010001100: z <= 10'b0000110000; // 4 * 12 = 48
            10'b0010001101: z <= 10'b0000110100; // 4 * 13 = 52
            10'b0010001110: z <= 10'b0000111000; // 4 * 14 = 56
            10'b0010001111: z <= 10'b0000111100; // 4 * 15 = 60
            10'b0010010000: z <= 10'b0001000000; // 4 * 16 = 64
            10'b0010010001: z <= 10'b0001000100; // 4 * 17 = 68
            10'b0010010010: z <= 10'b0001001000; // 4 * 18 = 72
            10'b0010010011: z <= 10'b0001001100; // 4 * 19 = 76
            10'b0010010100: z <= 10'b0001010000; // 4 * 20 = 80
            10'b0010010101: z <= 10'b0001010100; // 4 * 21 = 84
            10'b0010010110: z <= 10'b0001011000; // 4 * 22 = 88
            10'b0010010111: z <= 10'b0001011100; // 4 * 23 = 92
            10'b0010011000: z <= 10'b0001100000; // 4 * 24 = 96
            10'b0010011001: z <= 10'b0001100100; // 4 * 25 = 100
            10'b0010011010: z <= 10'b0001101000; // 4 * 26 = 104
            10'b0010011011: z <= 10'b0001101100; // 4 * 27 = 108
            10'b0010011100: z <= 10'b0001110000; // 4 * 28 = 112
            10'b0010011101: z <= 10'b0001110100; // 4 * 29 = 116
            10'b0010011110: z <= 10'b0001111000; // 4 * 30 = 120
            10'b0010011111: z <= 10'b0001111100; // 4 * 31 = 124
            10'b0010100000: z <= 10'b0000000000; // 5 * 0 = 0
            10'b0010100001: z <= 10'b0000000101; // 5 * 1 = 5
            10'b0010100010: z <= 10'b0000001010; // 5 * 2 = 10
            10'b0010100011: z <= 10'b0000001111; // 5 * 3 = 15
            10'b0010100100: z <= 10'b0000010100; // 5 * 4 = 20
            10'b0010100101: z <= 10'b0000011001; // 5 * 5 = 25
            10'b0010100110: z <= 10'b0000011110; // 5 * 6 = 30
            10'b0010100111: z <= 10'b0000100011; // 5 * 7 = 35
            10'b0010101000: z <= 10'b0000101000; // 5 * 8 = 40
            10'b0010101001: z <= 10'b0000101101; // 5 * 9 = 45
            10'b0010101010: z <= 10'b0000110010; // 5 * 10 = 50
            10'b0010101011: z <= 10'b0000110111; // 5 * 11 = 55
            10'b0010101100: z <= 10'b0000111100; // 5 * 12 = 60
            10'b0010101101: z <= 10'b0001000001; // 5 * 13 = 65
            10'b0010101110: z <= 10'b0001000110; // 5 * 14 = 70
            10'b0010101111: z <= 10'b0001001011; // 5 * 15 = 75
            10'b0010110000: z <= 10'b0001010000; // 5 * 16 = 80
            10'b0010110001: z <= 10'b0001010101; // 5 * 17 = 85
            10'b0010110010: z <= 10'b0001011010; // 5 * 18 = 90
            10'b0010110011: z <= 10'b0001011111; // 5 * 19 = 95
            10'b0010110100: z <= 10'b0001100100; // 5 * 20 = 100
            10'b0010110101: z <= 10'b0001101001; // 5 * 21 = 105
            10'b0010110110: z <= 10'b0001101110; // 5 * 22 = 110
            10'b0010110111: z <= 10'b0001110011; // 5 * 23 = 115
            10'b0010111000: z <= 10'b0001111000; // 5 * 24 = 120
            10'b0010111001: z <= 10'b0001111101; // 5 * 25 = 125
            10'b0010111010: z <= 10'b0010000010; // 5 * 26 = 130
            10'b0010111011: z <= 10'b0010000111; // 5 * 27 = 135
            10'b0010111100: z <= 10'b0010001100; // 5 * 28 = 140
            10'b0010111101: z <= 10'b0010010001; // 5 * 29 = 145
            10'b0010111110: z <= 10'b0010010110; // 5 * 30 = 150
            10'b0010111111: z <= 10'b0010011011; // 5 * 31 = 155
            10'b0011000000: z <= 10'b0000000000; // 6 * 0 = 0
            10'b0011000001: z <= 10'b0000000110; // 6 * 1 = 6
            10'b0011000010: z <= 10'b0000001100; // 6 * 2 = 12
            10'b0011000011: z <= 10'b0000010010; // 6 * 3 = 18
            10'b0011000100: z <= 10'b0000011000; // 6 * 4 = 24
            10'b0011000101: z <= 10'b0000011110; // 6 * 5 = 30
            10'b0011000110: z <= 10'b0000100100; // 6 * 6 = 36
            10'b0011000111: z <= 10'b0000101010; // 6 * 7 = 42
            10'b0011001000: z <= 10'b0000110000; // 6 * 8 = 48
            10'b0011001001: z <= 10'b0000110110; // 6 * 9 = 54
            10'b0011001010: z <= 10'b0000111100; // 6 * 10 = 60
            10'b0011001011: z <= 10'b0001000010; // 6 * 11 = 66
            10'b0011001100: z <= 10'b0001001000; // 6 * 12 = 72
            10'b0011001101: z <= 10'b0001001110; // 6 * 13 = 78
            10'b0011001110: z <= 10'b0001010100; // 6 * 14 = 84
            10'b0011001111: z <= 10'b0001011010; // 6 * 15 = 90
            10'b0011010000: z <= 10'b0001100000; // 6 * 16 = 96
            10'b0011010001: z <= 10'b0001100110; // 6 * 17 = 102
            10'b0011010010: z <= 10'b0001101100; // 6 * 18 = 108
            10'b0011010011: z <= 10'b0001110010; // 6 * 19 = 114
            10'b0011010100: z <= 10'b0001111000; // 6 * 20 = 120
            10'b0011010101: z <= 10'b0001111110; // 6 * 21 = 126
            10'b0011010110: z <= 10'b0010000100; // 6 * 22 = 132
            10'b0011010111: z <= 10'b0010001010; // 6 * 23 = 138
            10'b0011011000: z <= 10'b0010010000; // 6 * 24 = 144
            10'b0011011001: z <= 10'b0010010110; // 6 * 25 = 150
            10'b0011011010: z <= 10'b0010011100; // 6 * 26 = 156
            10'b0011011011: z <= 10'b0010100010; // 6 * 27 = 162
            10'b0011011100: z <= 10'b0010101000; // 6 * 28 = 168
            10'b0011011101: z <= 10'b0010101110; // 6 * 29 = 174
            10'b0011011110: z <= 10'b0010110100; // 6 * 30 = 180
            10'b0011011111: z <= 10'b0010111010; // 6 * 31 = 186
            10'b0011100000: z <= 10'b0000000000; // 7 * 0 = 0
            10'b0011100001: z <= 10'b0000000111; // 7 * 1 = 7
            10'b0011100010: z <= 10'b0000001110; // 7 * 2 = 14
            10'b0011100011: z <= 10'b0000010101; // 7 * 3 = 21
            10'b0011100100: z <= 10'b0000011100; // 7 * 4 = 28
            10'b0011100101: z <= 10'b0000100011; // 7 * 5 = 35
            10'b0011100110: z <= 10'b0000101010; // 7 * 6 = 42
            10'b0011100111: z <= 10'b0000110001; // 7 * 7 = 49
            10'b0011101000: z <= 10'b0000111000; // 7 * 8 = 56
            10'b0011101001: z <= 10'b0000111111; // 7 * 9 = 63
            10'b0011101010: z <= 10'b0001000110; // 7 * 10 = 70
            10'b0011101011: z <= 10'b0001001101; // 7 * 11 = 77
            10'b0011101100: z <= 10'b0001010100; // 7 * 12 = 84
            10'b0011101101: z <= 10'b0001011011; // 7 * 13 = 91
            10'b0011101110: z <= 10'b0001100010; // 7 * 14 = 98
            10'b0011101111: z <= 10'b0001101001; // 7 * 15 = 105
            10'b0011110000: z <= 10'b0001110000; // 7 * 16 = 112
            10'b0011110001: z <= 10'b0001110111; // 7 * 17 = 119
            10'b0011110010: z <= 10'b0001111110; // 7 * 18 = 126
            10'b0011110011: z <= 10'b0010000101; // 7 * 19 = 133
            10'b0011110100: z <= 10'b0010001100; // 7 * 20 = 140
            10'b0011110101: z <= 10'b0010010011; // 7 * 21 = 147
            10'b0011110110: z <= 10'b0010011010; // 7 * 22 = 154
            10'b0011110111: z <= 10'b0010100001; // 7 * 23 = 161
            10'b0011111000: z <= 10'b0010101000; // 7 * 24 = 168
            10'b0011111001: z <= 10'b0010101111; // 7 * 25 = 175
            10'b0011111010: z <= 10'b0010110110; // 7 * 26 = 182
            10'b0011111011: z <= 10'b0010111101; // 7 * 27 = 189
            10'b0011111100: z <= 10'b0011000100; // 7 * 28 = 196
            10'b0011111101: z <= 10'b0011001011; // 7 * 29 = 203
            10'b0011111110: z <= 10'b0011010010; // 7 * 30 = 210
            10'b0011111111: z <= 10'b0011011001; // 7 * 31 = 217
            10'b0100000000: z <= 10'b0000000000; // 8 * 0 = 0
            10'b0100000001: z <= 10'b0000001000; // 8 * 1 = 8
            10'b0100000010: z <= 10'b0000010000; // 8 * 2 = 16
            10'b0100000011: z <= 10'b0000011000; // 8 * 3 = 24
            10'b0100000100: z <= 10'b0000100000; // 8 * 4 = 32
            10'b0100000101: z <= 10'b0000101000; // 8 * 5 = 40
            10'b0100000110: z <= 10'b0000110000; // 8 * 6 = 48
            10'b0100000111: z <= 10'b0000111000; // 8 * 7 = 56
            10'b0100001000: z <= 10'b0001000000; // 8 * 8 = 64
            10'b0100001001: z <= 10'b0001001000; // 8 * 9 = 72
            10'b0100001010: z <= 10'b0001010000; // 8 * 10 = 80
            10'b0100001011: z <= 10'b0001011000; // 8 * 11 = 88
            10'b0100001100: z <= 10'b0001100000; // 8 * 12 = 96
            10'b0100001101: z <= 10'b0001101000; // 8 * 13 = 104
            10'b0100001110: z <= 10'b0001110000; // 8 * 14 = 112
            10'b0100001111: z <= 10'b0001111000; // 8 * 15 = 120
            10'b0100010000: z <= 10'b0010000000; // 8 * 16 = 128
            10'b0100010001: z <= 10'b0010001000; // 8 * 17 = 136
            10'b0100010010: z <= 10'b0010010000; // 8 * 18 = 144
            10'b0100010011: z <= 10'b0010011000; // 8 * 19 = 152
            10'b0100010100: z <= 10'b0010100000; // 8 * 20 = 160
            10'b0100010101: z <= 10'b0010101000; // 8 * 21 = 168
            10'b0100010110: z <= 10'b0010110000; // 8 * 22 = 176
            10'b0100010111: z <= 10'b0010111000; // 8 * 23 = 184
            10'b0100011000: z <= 10'b0011000000; // 8 * 24 = 192
            10'b0100011001: z <= 10'b0011001000; // 8 * 25 = 200
            10'b0100011010: z <= 10'b0011010000; // 8 * 26 = 208
            10'b0100011011: z <= 10'b0011011000; // 8 * 27 = 216
            10'b0100011100: z <= 10'b0011100000; // 8 * 28 = 224
            10'b0100011101: z <= 10'b0011101000; // 8 * 29 = 232
            10'b0100011110: z <= 10'b0011110000; // 8 * 30 = 240
            10'b0100011111: z <= 10'b0011111000; // 8 * 31 = 248
            10'b0100100000: z <= 10'b0000000000; // 9 * 0 = 0
            10'b0100100001: z <= 10'b0000001001; // 9 * 1 = 9
            10'b0100100010: z <= 10'b0000010010; // 9 * 2 = 18
            10'b0100100011: z <= 10'b0000011011; // 9 * 3 = 27
            10'b0100100100: z <= 10'b0000100100; // 9 * 4 = 36
            10'b0100100101: z <= 10'b0000101101; // 9 * 5 = 45
            10'b0100100110: z <= 10'b0000110110; // 9 * 6 = 54
            10'b0100100111: z <= 10'b0000111111; // 9 * 7 = 63
            10'b0100101000: z <= 10'b0001001000; // 9 * 8 = 72
            10'b0100101001: z <= 10'b0001010001; // 9 * 9 = 81
            10'b0100101010: z <= 10'b0001011010; // 9 * 10 = 90
            10'b0100101011: z <= 10'b0001100011; // 9 * 11 = 99
            10'b0100101100: z <= 10'b0001101100; // 9 * 12 = 108
            10'b0100101101: z <= 10'b0001110101; // 9 * 13 = 117
            10'b0100101110: z <= 10'b0001111110; // 9 * 14 = 126
            10'b0100101111: z <= 10'b0010000111; // 9 * 15 = 135
            10'b0100110000: z <= 10'b0010010000; // 9 * 16 = 144
            10'b0100110001: z <= 10'b0010011001; // 9 * 17 = 153
            10'b0100110010: z <= 10'b0010100010; // 9 * 18 = 162
            10'b0100110011: z <= 10'b0010101011; // 9 * 19 = 171
            10'b0100110100: z <= 10'b0010110100; // 9 * 20 = 180
            10'b0100110101: z <= 10'b0010111101; // 9 * 21 = 189
            10'b0100110110: z <= 10'b0011000110; // 9 * 22 = 198
            10'b0100110111: z <= 10'b0011001111; // 9 * 23 = 207
            10'b0100111000: z <= 10'b0011011000; // 9 * 24 = 216
            10'b0100111001: z <= 10'b0011100001; // 9 * 25 = 225
            10'b0100111010: z <= 10'b0011101010; // 9 * 26 = 234
            10'b0100111011: z <= 10'b0011110011; // 9 * 27 = 243
            10'b0100111100: z <= 10'b0011111100; // 9 * 28 = 252
            10'b0100111101: z <= 10'b0100000101; // 9 * 29 = 261
            10'b0100111110: z <= 10'b0100001110; // 9 * 30 = 270
            10'b0100111111: z <= 10'b0100010111; // 9 * 31 = 279
            10'b0101000000: z <= 10'b0000000000; // 10 * 0 = 0
            10'b0101000001: z <= 10'b0000001010; // 10 * 1 = 10
            10'b0101000010: z <= 10'b0000010100; // 10 * 2 = 20
            10'b0101000011: z <= 10'b0000011110; // 10 * 3 = 30
            10'b0101000100: z <= 10'b0000101000; // 10 * 4 = 40
            10'b0101000101: z <= 10'b0000110010; // 10 * 5 = 50
            10'b0101000110: z <= 10'b0000111100; // 10 * 6 = 60
            10'b0101000111: z <= 10'b0001000110; // 10 * 7 = 70
            10'b0101001000: z <= 10'b0001010000; // 10 * 8 = 80
            10'b0101001001: z <= 10'b0001011010; // 10 * 9 = 90
            10'b0101001010: z <= 10'b0001100100; // 10 * 10 = 100
            10'b0101001011: z <= 10'b0001101110; // 10 * 11 = 110
            10'b0101001100: z <= 10'b0001111000; // 10 * 12 = 120
            10'b0101001101: z <= 10'b0010000010; // 10 * 13 = 130
            10'b0101001110: z <= 10'b0010001100; // 10 * 14 = 140
            10'b0101001111: z <= 10'b0010010110; // 10 * 15 = 150
            10'b0101010000: z <= 10'b0010100000; // 10 * 16 = 160
            10'b0101010001: z <= 10'b0010101010; // 10 * 17 = 170
            10'b0101010010: z <= 10'b0010110100; // 10 * 18 = 180
            10'b0101010011: z <= 10'b0010111110; // 10 * 19 = 190
            10'b0101010100: z <= 10'b0011001000; // 10 * 20 = 200
            10'b0101010101: z <= 10'b0011010010; // 10 * 21 = 210
            10'b0101010110: z <= 10'b0011011100; // 10 * 22 = 220
            10'b0101010111: z <= 10'b0011100110; // 10 * 23 = 230
            10'b0101011000: z <= 10'b0011110000; // 10 * 24 = 240
            10'b0101011001: z <= 10'b0011111010; // 10 * 25 = 250
            10'b0101011010: z <= 10'b0100000100; // 10 * 26 = 260
            10'b0101011011: z <= 10'b0100001110; // 10 * 27 = 270
            10'b0101011100: z <= 10'b0100011000; // 10 * 28 = 280
            10'b0101011101: z <= 10'b0100100010; // 10 * 29 = 290
            10'b0101011110: z <= 10'b0100101100; // 10 * 30 = 300
            10'b0101011111: z <= 10'b0100110110; // 10 * 31 = 310
            10'b0101100000: z <= 10'b0000000000; // 11 * 0 = 0
            10'b0101100001: z <= 10'b0000001011; // 11 * 1 = 11
            10'b0101100010: z <= 10'b0000010110; // 11 * 2 = 22
            10'b0101100011: z <= 10'b0000100001; // 11 * 3 = 33
            10'b0101100100: z <= 10'b0000101100; // 11 * 4 = 44
            10'b0101100101: z <= 10'b0000110111; // 11 * 5 = 55
            10'b0101100110: z <= 10'b0001000010; // 11 * 6 = 66
            10'b0101100111: z <= 10'b0001001101; // 11 * 7 = 77
            10'b0101101000: z <= 10'b0001011000; // 11 * 8 = 88
            10'b0101101001: z <= 10'b0001100011; // 11 * 9 = 99
            10'b0101101010: z <= 10'b0001101110; // 11 * 10 = 110
            10'b0101101011: z <= 10'b0001111001; // 11 * 11 = 121
            10'b0101101100: z <= 10'b0010000100; // 11 * 12 = 132
            10'b0101101101: z <= 10'b0010001111; // 11 * 13 = 143
            10'b0101101110: z <= 10'b0010011010; // 11 * 14 = 154
            10'b0101101111: z <= 10'b0010100101; // 11 * 15 = 165
            10'b0101110000: z <= 10'b0010110000; // 11 * 16 = 176
            10'b0101110001: z <= 10'b0010111011; // 11 * 17 = 187
            10'b0101110010: z <= 10'b0011000110; // 11 * 18 = 198
            10'b0101110011: z <= 10'b0011010001; // 11 * 19 = 209
            10'b0101110100: z <= 10'b0011011100; // 11 * 20 = 220
            10'b0101110101: z <= 10'b0011100111; // 11 * 21 = 231
            10'b0101110110: z <= 10'b0011110010; // 11 * 22 = 242
            10'b0101110111: z <= 10'b0011111101; // 11 * 23 = 253
            10'b0101111000: z <= 10'b0100001000; // 11 * 24 = 264
            10'b0101111001: z <= 10'b0100010011; // 11 * 25 = 275
            10'b0101111010: z <= 10'b0100011110; // 11 * 26 = 286
            10'b0101111011: z <= 10'b0100101001; // 11 * 27 = 297
            10'b0101111100: z <= 10'b0100110100; // 11 * 28 = 308
            10'b0101111101: z <= 10'b0100111111; // 11 * 29 = 319
            10'b0101111110: z <= 10'b0101001010; // 11 * 30 = 330
            10'b0101111111: z <= 10'b0101010101; // 11 * 31 = 341
            10'b0110000000: z <= 10'b0000000000; // 12 * 0 = 0
            10'b0110000001: z <= 10'b0000001100; // 12 * 1 = 12
            10'b0110000010: z <= 10'b0000011000; // 12 * 2 = 24
            10'b0110000011: z <= 10'b0000100100; // 12 * 3 = 36
            10'b0110000100: z <= 10'b0000110000; // 12 * 4 = 48
            10'b0110000101: z <= 10'b0000111100; // 12 * 5 = 60
            10'b0110000110: z <= 10'b0001001000; // 12 * 6 = 72
            10'b0110000111: z <= 10'b0001010100; // 12 * 7 = 84
            10'b0110001000: z <= 10'b0001100000; // 12 * 8 = 96
            10'b0110001001: z <= 10'b0001101100; // 12 * 9 = 108
            10'b0110001010: z <= 10'b0001111000; // 12 * 10 = 120
            10'b0110001011: z <= 10'b0010000100; // 12 * 11 = 132
            10'b0110001100: z <= 10'b0010010000; // 12 * 12 = 144
            10'b0110001101: z <= 10'b0010011100; // 12 * 13 = 156
            10'b0110001110: z <= 10'b0010101000; // 12 * 14 = 168
            10'b0110001111: z <= 10'b0010110100; // 12 * 15 = 180
            10'b0110010000: z <= 10'b0011000000; // 12 * 16 = 192
            10'b0110010001: z <= 10'b0011001100; // 12 * 17 = 204
            10'b0110010010: z <= 10'b0011011000; // 12 * 18 = 216
            10'b0110010011: z <= 10'b0011100100; // 12 * 19 = 228
            10'b0110010100: z <= 10'b0011110000; // 12 * 20 = 240
            10'b0110010101: z <= 10'b0011111100; // 12 * 21 = 252
            10'b0110010110: z <= 10'b0100001000; // 12 * 22 = 264
            10'b0110010111: z <= 10'b0100010100; // 12 * 23 = 276
            10'b0110011000: z <= 10'b0100100000; // 12 * 24 = 288
            10'b0110011001: z <= 10'b0100101100; // 12 * 25 = 300
            10'b0110011010: z <= 10'b0100111000; // 12 * 26 = 312
            10'b0110011011: z <= 10'b0101000100; // 12 * 27 = 324
            10'b0110011100: z <= 10'b0101010000; // 12 * 28 = 336
            10'b0110011101: z <= 10'b0101011100; // 12 * 29 = 348
            10'b0110011110: z <= 10'b0101101000; // 12 * 30 = 360
            10'b0110011111: z <= 10'b0101110100; // 12 * 31 = 372
            10'b0110100000: z <= 10'b0000000000; // 13 * 0 = 0
            10'b0110100001: z <= 10'b0000001101; // 13 * 1 = 13
            10'b0110100010: z <= 10'b0000011010; // 13 * 2 = 26
            10'b0110100011: z <= 10'b0000100111; // 13 * 3 = 39
            10'b0110100100: z <= 10'b0000110100; // 13 * 4 = 52
            10'b0110100101: z <= 10'b0001000001; // 13 * 5 = 65
            10'b0110100110: z <= 10'b0001001110; // 13 * 6 = 78
            10'b0110100111: z <= 10'b0001011011; // 13 * 7 = 91
            10'b0110101000: z <= 10'b0001101000; // 13 * 8 = 104
            10'b0110101001: z <= 10'b0001110101; // 13 * 9 = 117
            10'b0110101010: z <= 10'b0010000010; // 13 * 10 = 130
            10'b0110101011: z <= 10'b0010001111; // 13 * 11 = 143
            10'b0110101100: z <= 10'b0010011100; // 13 * 12 = 156
            10'b0110101101: z <= 10'b0010101001; // 13 * 13 = 169
            10'b0110101110: z <= 10'b0010110110; // 13 * 14 = 182
            10'b0110101111: z <= 10'b0011000011; // 13 * 15 = 195
            10'b0110110000: z <= 10'b0011010000; // 13 * 16 = 208
            10'b0110110001: z <= 10'b0011011101; // 13 * 17 = 221
            10'b0110110010: z <= 10'b0011101010; // 13 * 18 = 234
            10'b0110110011: z <= 10'b0011110111; // 13 * 19 = 247
            10'b0110110100: z <= 10'b0100000100; // 13 * 20 = 260
            10'b0110110101: z <= 10'b0100010001; // 13 * 21 = 273
            10'b0110110110: z <= 10'b0100011110; // 13 * 22 = 286
            10'b0110110111: z <= 10'b0100101011; // 13 * 23 = 299
            10'b0110111000: z <= 10'b0100111000; // 13 * 24 = 312
            10'b0110111001: z <= 10'b0101000101; // 13 * 25 = 325
            10'b0110111010: z <= 10'b0101010010; // 13 * 26 = 338
            10'b0110111011: z <= 10'b0101011111; // 13 * 27 = 351
            10'b0110111100: z <= 10'b0101101100; // 13 * 28 = 364
            10'b0110111101: z <= 10'b0101111001; // 13 * 29 = 377
            10'b0110111110: z <= 10'b0110000110; // 13 * 30 = 390
            10'b0110111111: z <= 10'b0110010011; // 13 * 31 = 403
            10'b0111000000: z <= 10'b0000000000; // 14 * 0 = 0
            10'b0111000001: z <= 10'b0000001110; // 14 * 1 = 14
            10'b0111000010: z <= 10'b0000011100; // 14 * 2 = 28
            10'b0111000011: z <= 10'b0000101010; // 14 * 3 = 42
            10'b0111000100: z <= 10'b0000111000; // 14 * 4 = 56
            10'b0111000101: z <= 10'b0001000110; // 14 * 5 = 70
            10'b0111000110: z <= 10'b0001010100; // 14 * 6 = 84
            10'b0111000111: z <= 10'b0001100010; // 14 * 7 = 98
            10'b0111001000: z <= 10'b0001110000; // 14 * 8 = 112
            10'b0111001001: z <= 10'b0001111110; // 14 * 9 = 126
            10'b0111001010: z <= 10'b0010001100; // 14 * 10 = 140
            10'b0111001011: z <= 10'b0010011010; // 14 * 11 = 154
            10'b0111001100: z <= 10'b0010101000; // 14 * 12 = 168
            10'b0111001101: z <= 10'b0010110110; // 14 * 13 = 182
            10'b0111001110: z <= 10'b0011000100; // 14 * 14 = 196
            10'b0111001111: z <= 10'b0011010010; // 14 * 15 = 210
            10'b0111010000: z <= 10'b0011100000; // 14 * 16 = 224
            10'b0111010001: z <= 10'b0011101110; // 14 * 17 = 238
            10'b0111010010: z <= 10'b0011111100; // 14 * 18 = 252
            10'b0111010011: z <= 10'b0100001010; // 14 * 19 = 266
            10'b0111010100: z <= 10'b0100011000; // 14 * 20 = 280
            10'b0111010101: z <= 10'b0100100110; // 14 * 21 = 294
            10'b0111010110: z <= 10'b0100110100; // 14 * 22 = 308
            10'b0111010111: z <= 10'b0101000010; // 14 * 23 = 322
            10'b0111011000: z <= 10'b0101010000; // 14 * 24 = 336
            10'b0111011001: z <= 10'b0101011110; // 14 * 25 = 350
            10'b0111011010: z <= 10'b0101101100; // 14 * 26 = 364
            10'b0111011011: z <= 10'b0101111010; // 14 * 27 = 378
            10'b0111011100: z <= 10'b0110001000; // 14 * 28 = 392
            10'b0111011101: z <= 10'b0110010110; // 14 * 29 = 406
            10'b0111011110: z <= 10'b0110100100; // 14 * 30 = 420
            10'b0111011111: z <= 10'b0110110010; // 14 * 31 = 434
            10'b0111100000: z <= 10'b0000000000; // 15 * 0 = 0
            10'b0111100001: z <= 10'b0000001111; // 15 * 1 = 15
            10'b0111100010: z <= 10'b0000011110; // 15 * 2 = 30
            10'b0111100011: z <= 10'b0000101101; // 15 * 3 = 45
            10'b0111100100: z <= 10'b0000111100; // 15 * 4 = 60
            10'b0111100101: z <= 10'b0001001011; // 15 * 5 = 75
            10'b0111100110: z <= 10'b0001011010; // 15 * 6 = 90
            10'b0111100111: z <= 10'b0001101001; // 15 * 7 = 105
            10'b0111101000: z <= 10'b0001111000; // 15 * 8 = 120
            10'b0111101001: z <= 10'b0010000111; // 15 * 9 = 135
            10'b0111101010: z <= 10'b0010010110; // 15 * 10 = 150
            10'b0111101011: z <= 10'b0010100101; // 15 * 11 = 165
            10'b0111101100: z <= 10'b0010110100; // 15 * 12 = 180
            10'b0111101101: z <= 10'b0011000011; // 15 * 13 = 195
            10'b0111101110: z <= 10'b0011010010; // 15 * 14 = 210
            10'b0111101111: z <= 10'b0011100001; // 15 * 15 = 225
            10'b0111110000: z <= 10'b0011110000; // 15 * 16 = 240
            10'b0111110001: z <= 10'b0011111111; // 15 * 17 = 255
            10'b0111110010: z <= 10'b0100001110; // 15 * 18 = 270
            10'b0111110011: z <= 10'b0100011101; // 15 * 19 = 285
            10'b0111110100: z <= 10'b0100101100; // 15 * 20 = 300
            10'b0111110101: z <= 10'b0100111011; // 15 * 21 = 315
            10'b0111110110: z <= 10'b0101001010; // 15 * 22 = 330
            10'b0111110111: z <= 10'b0101011001; // 15 * 23 = 345
            10'b0111111000: z <= 10'b0101101000; // 15 * 24 = 360
            10'b0111111001: z <= 10'b0101110111; // 15 * 25 = 375
            10'b0111111010: z <= 10'b0110000110; // 15 * 26 = 390
            10'b0111111011: z <= 10'b0110010101; // 15 * 27 = 405
            10'b0111111100: z <= 10'b0110100100; // 15 * 28 = 420
            10'b0111111101: z <= 10'b0110110011; // 15 * 29 = 435
            10'b0111111110: z <= 10'b0111000010; // 15 * 30 = 450
            10'b0111111111: z <= 10'b0111010001; // 15 * 31 = 465
            10'b1000000000: z <= 10'b0000000000; // 16 * 0 = 0
            10'b1000000001: z <= 10'b0000010000; // 16 * 1 = 16
            10'b1000000010: z <= 10'b0000100000; // 16 * 2 = 32
            10'b1000000011: z <= 10'b0000110000; // 16 * 3 = 48
            10'b1000000100: z <= 10'b0001000000; // 16 * 4 = 64
            10'b1000000101: z <= 10'b0001010000; // 16 * 5 = 80
            10'b1000000110: z <= 10'b0001100000; // 16 * 6 = 96
            10'b1000000111: z <= 10'b0001110000; // 16 * 7 = 112
            10'b1000001000: z <= 10'b0010000000; // 16 * 8 = 128
            10'b1000001001: z <= 10'b0010010000; // 16 * 9 = 144
            10'b1000001010: z <= 10'b0010100000; // 16 * 10 = 160
            10'b1000001011: z <= 10'b0010110000; // 16 * 11 = 176
            10'b1000001100: z <= 10'b0011000000; // 16 * 12 = 192
            10'b1000001101: z <= 10'b0011010000; // 16 * 13 = 208
            10'b1000001110: z <= 10'b0011100000; // 16 * 14 = 224
            10'b1000001111: z <= 10'b0011110000; // 16 * 15 = 240
            10'b1000010000: z <= 10'b0100000000; // 16 * 16 = 256
            10'b1000010001: z <= 10'b0100010000; // 16 * 17 = 272
            10'b1000010010: z <= 10'b0100100000; // 16 * 18 = 288
            10'b1000010011: z <= 10'b0100110000; // 16 * 19 = 304
            10'b1000010100: z <= 10'b0101000000; // 16 * 20 = 320
            10'b1000010101: z <= 10'b0101010000; // 16 * 21 = 336
            10'b1000010110: z <= 10'b0101100000; // 16 * 22 = 352
            10'b1000010111: z <= 10'b0101110000; // 16 * 23 = 368
            10'b1000011000: z <= 10'b0110000000; // 16 * 24 = 384
            10'b1000011001: z <= 10'b0110010000; // 16 * 25 = 400
            10'b1000011010: z <= 10'b0110100000; // 16 * 26 = 416
            10'b1000011011: z <= 10'b0110110000; // 16 * 27 = 432
            10'b1000011100: z <= 10'b0111000000; // 16 * 28 = 448
            10'b1000011101: z <= 10'b0111010000; // 16 * 29 = 464
            10'b1000011110: z <= 10'b0111100000; // 16 * 30 = 480
            10'b1000011111: z <= 10'b0111110000; // 16 * 31 = 496
            10'b1000100000: z <= 10'b0000000000; // 17 * 0 = 0
            10'b1000100001: z <= 10'b0000010001; // 17 * 1 = 17
            10'b1000100010: z <= 10'b0000100010; // 17 * 2 = 34
            10'b1000100011: z <= 10'b0000110011; // 17 * 3 = 51
            10'b1000100100: z <= 10'b0001000100; // 17 * 4 = 68
            10'b1000100101: z <= 10'b0001010101; // 17 * 5 = 85
            10'b1000100110: z <= 10'b0001100110; // 17 * 6 = 102
            10'b1000100111: z <= 10'b0001110111; // 17 * 7 = 119
            10'b1000101000: z <= 10'b0010001000; // 17 * 8 = 136
            10'b1000101001: z <= 10'b0010011001; // 17 * 9 = 153
            10'b1000101010: z <= 10'b0010101010; // 17 * 10 = 170
            10'b1000101011: z <= 10'b0010111011; // 17 * 11 = 187
            10'b1000101100: z <= 10'b0011001100; // 17 * 12 = 204
            10'b1000101101: z <= 10'b0011011101; // 17 * 13 = 221
            10'b1000101110: z <= 10'b0011101110; // 17 * 14 = 238
            10'b1000101111: z <= 10'b0011111111; // 17 * 15 = 255
            10'b1000110000: z <= 10'b0100010000; // 17 * 16 = 272
            10'b1000110001: z <= 10'b0100100001; // 17 * 17 = 289
            10'b1000110010: z <= 10'b0100110010; // 17 * 18 = 306
            10'b1000110011: z <= 10'b0101000011; // 17 * 19 = 323
            10'b1000110100: z <= 10'b0101010100; // 17 * 20 = 340
            10'b1000110101: z <= 10'b0101100101; // 17 * 21 = 357
            10'b1000110110: z <= 10'b0101110110; // 17 * 22 = 374
            10'b1000110111: z <= 10'b0110000111; // 17 * 23 = 391
            10'b1000111000: z <= 10'b0110011000; // 17 * 24 = 408
            10'b1000111001: z <= 10'b0110101001; // 17 * 25 = 425
            10'b1000111010: z <= 10'b0110111010; // 17 * 26 = 442
            10'b1000111011: z <= 10'b0111001011; // 17 * 27 = 459
            10'b1000111100: z <= 10'b0111011100; // 17 * 28 = 476
            10'b1000111101: z <= 10'b0111101101; // 17 * 29 = 493
            10'b1000111110: z <= 10'b0111111110; // 17 * 30 = 510
            10'b1000111111: z <= 10'b1000001111; // 17 * 31 = 527
            10'b1001000000: z <= 10'b0000000000; // 18 * 0 = 0
            10'b1001000001: z <= 10'b0000010010; // 18 * 1 = 18
            10'b1001000010: z <= 10'b0000100100; // 18 * 2 = 36
            10'b1001000011: z <= 10'b0000110110; // 18 * 3 = 54
            10'b1001000100: z <= 10'b0001001000; // 18 * 4 = 72
            10'b1001000101: z <= 10'b0001011010; // 18 * 5 = 90
            10'b1001000110: z <= 10'b0001101100; // 18 * 6 = 108
            10'b1001000111: z <= 10'b0001111110; // 18 * 7 = 126
            10'b1001001000: z <= 10'b0010010000; // 18 * 8 = 144
            10'b1001001001: z <= 10'b0010100010; // 18 * 9 = 162
            10'b1001001010: z <= 10'b0010110100; // 18 * 10 = 180
            10'b1001001011: z <= 10'b0011000110; // 18 * 11 = 198
            10'b1001001100: z <= 10'b0011011000; // 18 * 12 = 216
            10'b1001001101: z <= 10'b0011101010; // 18 * 13 = 234
            10'b1001001110: z <= 10'b0011111100; // 18 * 14 = 252
            10'b1001001111: z <= 10'b0100001110; // 18 * 15 = 270
            10'b1001010000: z <= 10'b0100100000; // 18 * 16 = 288
            10'b1001010001: z <= 10'b0100110010; // 18 * 17 = 306
            10'b1001010010: z <= 10'b0101000100; // 18 * 18 = 324
            10'b1001010011: z <= 10'b0101010110; // 18 * 19 = 342
            10'b1001010100: z <= 10'b0101101000; // 18 * 20 = 360
            10'b1001010101: z <= 10'b0101111010; // 18 * 21 = 378
            10'b1001010110: z <= 10'b0110001100; // 18 * 22 = 396
            10'b1001010111: z <= 10'b0110011110; // 18 * 23 = 414
            10'b1001011000: z <= 10'b0110110000; // 18 * 24 = 432
            10'b1001011001: z <= 10'b0111000010; // 18 * 25 = 450
            10'b1001011010: z <= 10'b0111010100; // 18 * 26 = 468
            10'b1001011011: z <= 10'b0111100110; // 18 * 27 = 486
            10'b1001011100: z <= 10'b0111111000; // 18 * 28 = 504
            10'b1001011101: z <= 10'b1000001010; // 18 * 29 = 522
            10'b1001011110: z <= 10'b1000011100; // 18 * 30 = 540
            10'b1001011111: z <= 10'b1000101110; // 18 * 31 = 558
            10'b1001100000: z <= 10'b0000000000; // 19 * 0 = 0
            10'b1001100001: z <= 10'b0000010011; // 19 * 1 = 19
            10'b1001100010: z <= 10'b0000100110; // 19 * 2 = 38
            10'b1001100011: z <= 10'b0000111001; // 19 * 3 = 57
            10'b1001100100: z <= 10'b0001001100; // 19 * 4 = 76
            10'b1001100101: z <= 10'b0001011111; // 19 * 5 = 95
            10'b1001100110: z <= 10'b0001110010; // 19 * 6 = 114
            10'b1001100111: z <= 10'b0010000101; // 19 * 7 = 133
            10'b1001101000: z <= 10'b0010011000; // 19 * 8 = 152
            10'b1001101001: z <= 10'b0010101011; // 19 * 9 = 171
            10'b1001101010: z <= 10'b0010111110; // 19 * 10 = 190
            10'b1001101011: z <= 10'b0011010001; // 19 * 11 = 209
            10'b1001101100: z <= 10'b0011100100; // 19 * 12 = 228
            10'b1001101101: z <= 10'b0011110111; // 19 * 13 = 247
            10'b1001101110: z <= 10'b0100001010; // 19 * 14 = 266
            10'b1001101111: z <= 10'b0100011101; // 19 * 15 = 285
            10'b1001110000: z <= 10'b0100110000; // 19 * 16 = 304
            10'b1001110001: z <= 10'b0101000011; // 19 * 17 = 323
            10'b1001110010: z <= 10'b0101010110; // 19 * 18 = 342
            10'b1001110011: z <= 10'b0101101001; // 19 * 19 = 361
            10'b1001110100: z <= 10'b0101111100; // 19 * 20 = 380
            10'b1001110101: z <= 10'b0110001111; // 19 * 21 = 399
            10'b1001110110: z <= 10'b0110100010; // 19 * 22 = 418
            10'b1001110111: z <= 10'b0110110101; // 19 * 23 = 437
            10'b1001111000: z <= 10'b0111001000; // 19 * 24 = 456
            10'b1001111001: z <= 10'b0111011011; // 19 * 25 = 475
            10'b1001111010: z <= 10'b0111101110; // 19 * 26 = 494
            10'b1001111011: z <= 10'b1000000001; // 19 * 27 = 513
            10'b1001111100: z <= 10'b1000010100; // 19 * 28 = 532
            10'b1001111101: z <= 10'b1000100111; // 19 * 29 = 551
            10'b1001111110: z <= 10'b1000111010; // 19 * 30 = 570
            10'b1001111111: z <= 10'b1001001101; // 19 * 31 = 589
            10'b1010000000: z <= 10'b0000000000; // 20 * 0 = 0
            10'b1010000001: z <= 10'b0000010100; // 20 * 1 = 20
            10'b1010000010: z <= 10'b0000101000; // 20 * 2 = 40
            10'b1010000011: z <= 10'b0000111100; // 20 * 3 = 60
            10'b1010000100: z <= 10'b0001010000; // 20 * 4 = 80
            10'b1010000101: z <= 10'b0001100100; // 20 * 5 = 100
            10'b1010000110: z <= 10'b0001111000; // 20 * 6 = 120
            10'b1010000111: z <= 10'b0010001100; // 20 * 7 = 140
            10'b1010001000: z <= 10'b0010100000; // 20 * 8 = 160
            10'b1010001001: z <= 10'b0010110100; // 20 * 9 = 180
            10'b1010001010: z <= 10'b0011001000; // 20 * 10 = 200
            10'b1010001011: z <= 10'b0011011100; // 20 * 11 = 220
            10'b1010001100: z <= 10'b0011110000; // 20 * 12 = 240
            10'b1010001101: z <= 10'b0100000100; // 20 * 13 = 260
            10'b1010001110: z <= 10'b0100011000; // 20 * 14 = 280
            10'b1010001111: z <= 10'b0100101100; // 20 * 15 = 300
            10'b1010010000: z <= 10'b0101000000; // 20 * 16 = 320
            10'b1010010001: z <= 10'b0101010100; // 20 * 17 = 340
            10'b1010010010: z <= 10'b0101101000; // 20 * 18 = 360
            10'b1010010011: z <= 10'b0101111100; // 20 * 19 = 380
            10'b1010010100: z <= 10'b0110010000; // 20 * 20 = 400
            10'b1010010101: z <= 10'b0110100100; // 20 * 21 = 420
            10'b1010010110: z <= 10'b0110111000; // 20 * 22 = 440
            10'b1010010111: z <= 10'b0111001100; // 20 * 23 = 460
            10'b1010011000: z <= 10'b0111100000; // 20 * 24 = 480
            10'b1010011001: z <= 10'b0111110100; // 20 * 25 = 500
            10'b1010011010: z <= 10'b1000001000; // 20 * 26 = 520
            10'b1010011011: z <= 10'b1000011100; // 20 * 27 = 540
            10'b1010011100: z <= 10'b1000110000; // 20 * 28 = 560
            10'b1010011101: z <= 10'b1001000100; // 20 * 29 = 580
            10'b1010011110: z <= 10'b1001011000; // 20 * 30 = 600
            10'b1010011111: z <= 10'b1001101100; // 20 * 31 = 620
            10'b1010100000: z <= 10'b0000000000; // 21 * 0 = 0
            10'b1010100001: z <= 10'b0000010101; // 21 * 1 = 21
            10'b1010100010: z <= 10'b0000101010; // 21 * 2 = 42
            10'b1010100011: z <= 10'b0000111111; // 21 * 3 = 63
            10'b1010100100: z <= 10'b0001010100; // 21 * 4 = 84
            10'b1010100101: z <= 10'b0001101001; // 21 * 5 = 105
            10'b1010100110: z <= 10'b0001111110; // 21 * 6 = 126
            10'b1010100111: z <= 10'b0010010011; // 21 * 7 = 147
            10'b1010101000: z <= 10'b0010101000; // 21 * 8 = 168
            10'b1010101001: z <= 10'b0010111101; // 21 * 9 = 189
            10'b1010101010: z <= 10'b0011010010; // 21 * 10 = 210
            10'b1010101011: z <= 10'b0011100111; // 21 * 11 = 231
            10'b1010101100: z <= 10'b0011111100; // 21 * 12 = 252
            10'b1010101101: z <= 10'b0100010001; // 21 * 13 = 273
            10'b1010101110: z <= 10'b0100100110; // 21 * 14 = 294
            10'b1010101111: z <= 10'b0100111011; // 21 * 15 = 315
            10'b1010110000: z <= 10'b0101010000; // 21 * 16 = 336
            10'b1010110001: z <= 10'b0101100101; // 21 * 17 = 357
            10'b1010110010: z <= 10'b0101111010; // 21 * 18 = 378
            10'b1010110011: z <= 10'b0110001111; // 21 * 19 = 399
            10'b1010110100: z <= 10'b0110100100; // 21 * 20 = 420
            10'b1010110101: z <= 10'b0110111001; // 21 * 21 = 441
            10'b1010110110: z <= 10'b0111001110; // 21 * 22 = 462
            10'b1010110111: z <= 10'b0111100011; // 21 * 23 = 483
            10'b1010111000: z <= 10'b0111111000; // 21 * 24 = 504
            10'b1010111001: z <= 10'b1000001101; // 21 * 25 = 525
            10'b1010111010: z <= 10'b1000100010; // 21 * 26 = 546
            10'b1010111011: z <= 10'b1000110111; // 21 * 27 = 567
            10'b1010111100: z <= 10'b1001001100; // 21 * 28 = 588
            10'b1010111101: z <= 10'b1001100001; // 21 * 29 = 609
            10'b1010111110: z <= 10'b1001110110; // 21 * 30 = 630
            10'b1010111111: z <= 10'b1010001011; // 21 * 31 = 651
            10'b1011000000: z <= 10'b0000000000; // 22 * 0 = 0
            10'b1011000001: z <= 10'b0000010110; // 22 * 1 = 22
            10'b1011000010: z <= 10'b0000101100; // 22 * 2 = 44
            10'b1011000011: z <= 10'b0001000010; // 22 * 3 = 66
            10'b1011000100: z <= 10'b0001011000; // 22 * 4 = 88
            10'b1011000101: z <= 10'b0001101110; // 22 * 5 = 110
            10'b1011000110: z <= 10'b0010000100; // 22 * 6 = 132
            10'b1011000111: z <= 10'b0010011010; // 22 * 7 = 154
            10'b1011001000: z <= 10'b0010110000; // 22 * 8 = 176
            10'b1011001001: z <= 10'b0011000110; // 22 * 9 = 198
            10'b1011001010: z <= 10'b0011011100; // 22 * 10 = 220
            10'b1011001011: z <= 10'b0011110010; // 22 * 11 = 242
            10'b1011001100: z <= 10'b0100001000; // 22 * 12 = 264
            10'b1011001101: z <= 10'b0100011110; // 22 * 13 = 286
            10'b1011001110: z <= 10'b0100110100; // 22 * 14 = 308
            10'b1011001111: z <= 10'b0101001010; // 22 * 15 = 330
            10'b1011010000: z <= 10'b0101100000; // 22 * 16 = 352
            10'b1011010001: z <= 10'b0101110110; // 22 * 17 = 374
            10'b1011010010: z <= 10'b0110001100; // 22 * 18 = 396
            10'b1011010011: z <= 10'b0110100010; // 22 * 19 = 418
            10'b1011010100: z <= 10'b0110111000; // 22 * 20 = 440
            10'b1011010101: z <= 10'b0111001110; // 22 * 21 = 462
            10'b1011010110: z <= 10'b0111100100; // 22 * 22 = 484
            10'b1011010111: z <= 10'b0111111010; // 22 * 23 = 506
            10'b1011011000: z <= 10'b1000010000; // 22 * 24 = 528
            10'b1011011001: z <= 10'b1000100110; // 22 * 25 = 550
            10'b1011011010: z <= 10'b1000111100; // 22 * 26 = 572
            10'b1011011011: z <= 10'b1001010010; // 22 * 27 = 594
            10'b1011011100: z <= 10'b1001101000; // 22 * 28 = 616
            10'b1011011101: z <= 10'b1001111110; // 22 * 29 = 638
            10'b1011011110: z <= 10'b1010010100; // 22 * 30 = 660
            10'b1011011111: z <= 10'b1010101010; // 22 * 31 = 682
            10'b1011100000: z <= 10'b0000000000; // 23 * 0 = 0
            10'b1011100001: z <= 10'b0000010111; // 23 * 1 = 23
            10'b1011100010: z <= 10'b0000101110; // 23 * 2 = 46
            10'b1011100011: z <= 10'b0001000101; // 23 * 3 = 69
            10'b1011100100: z <= 10'b0001011100; // 23 * 4 = 92
            10'b1011100101: z <= 10'b0001110011; // 23 * 5 = 115
            10'b1011100110: z <= 10'b0010001010; // 23 * 6 = 138
            10'b1011100111: z <= 10'b0010100001; // 23 * 7 = 161
            10'b1011101000: z <= 10'b0010111000; // 23 * 8 = 184
            10'b1011101001: z <= 10'b0011001111; // 23 * 9 = 207
            10'b1011101010: z <= 10'b0011100110; // 23 * 10 = 230
            10'b1011101011: z <= 10'b0011111101; // 23 * 11 = 253
            10'b1011101100: z <= 10'b0100010100; // 23 * 12 = 276
            10'b1011101101: z <= 10'b0100101011; // 23 * 13 = 299
            10'b1011101110: z <= 10'b0101000010; // 23 * 14 = 322
            10'b1011101111: z <= 10'b0101011001; // 23 * 15 = 345
            10'b1011110000: z <= 10'b0101110000; // 23 * 16 = 368
            10'b1011110001: z <= 10'b0110000111; // 23 * 17 = 391
            10'b1011110010: z <= 10'b0110011110; // 23 * 18 = 414
            10'b1011110011: z <= 10'b0110110101; // 23 * 19 = 437
            10'b1011110100: z <= 10'b0111001100; // 23 * 20 = 460
            10'b1011110101: z <= 10'b0111100011; // 23 * 21 = 483
            10'b1011110110: z <= 10'b0111111010; // 23 * 22 = 506
            10'b1011110111: z <= 10'b1000010001; // 23 * 23 = 529
            10'b1011111000: z <= 10'b1000101000; // 23 * 24 = 552
            10'b1011111001: z <= 10'b1000111111; // 23 * 25 = 575
            10'b1011111010: z <= 10'b1001010110; // 23 * 26 = 598
            10'b1011111011: z <= 10'b1001101101; // 23 * 27 = 621
            10'b1011111100: z <= 10'b1010000100; // 23 * 28 = 644
            10'b1011111101: z <= 10'b1010011011; // 23 * 29 = 667
            10'b1011111110: z <= 10'b1010110010; // 23 * 30 = 690
            10'b1011111111: z <= 10'b1011001001; // 23 * 31 = 713
            10'b1100000000: z <= 10'b0000000000; // 24 * 0 = 0
            10'b1100000001: z <= 10'b0000011000; // 24 * 1 = 24
            10'b1100000010: z <= 10'b0000110000; // 24 * 2 = 48
            10'b1100000011: z <= 10'b0001001000; // 24 * 3 = 72
            10'b1100000100: z <= 10'b0001100000; // 24 * 4 = 96
            10'b1100000101: z <= 10'b0001111000; // 24 * 5 = 120
            10'b1100000110: z <= 10'b0010010000; // 24 * 6 = 144
            10'b1100000111: z <= 10'b0010101000; // 24 * 7 = 168
            10'b1100001000: z <= 10'b0011000000; // 24 * 8 = 192
            10'b1100001001: z <= 10'b0011011000; // 24 * 9 = 216
            10'b1100001010: z <= 10'b0011110000; // 24 * 10 = 240
            10'b1100001011: z <= 10'b0100001000; // 24 * 11 = 264
            10'b1100001100: z <= 10'b0100100000; // 24 * 12 = 288
            10'b1100001101: z <= 10'b0100111000; // 24 * 13 = 312
            10'b1100001110: z <= 10'b0101010000; // 24 * 14 = 336
            10'b1100001111: z <= 10'b0101101000; // 24 * 15 = 360
            10'b1100010000: z <= 10'b0110000000; // 24 * 16 = 384
            10'b1100010001: z <= 10'b0110011000; // 24 * 17 = 408
            10'b1100010010: z <= 10'b0110110000; // 24 * 18 = 432
            10'b1100010011: z <= 10'b0111001000; // 24 * 19 = 456
            10'b1100010100: z <= 10'b0111100000; // 24 * 20 = 480
            10'b1100010101: z <= 10'b0111111000; // 24 * 21 = 504
            10'b1100010110: z <= 10'b1000010000; // 24 * 22 = 528
            10'b1100010111: z <= 10'b1000101000; // 24 * 23 = 552
            10'b1100011000: z <= 10'b1001000000; // 24 * 24 = 576
            10'b1100011001: z <= 10'b1001011000; // 24 * 25 = 600
            10'b1100011010: z <= 10'b1001110000; // 24 * 26 = 624
            10'b1100011011: z <= 10'b1010001000; // 24 * 27 = 648
            10'b1100011100: z <= 10'b1010100000; // 24 * 28 = 672
            10'b1100011101: z <= 10'b1010111000; // 24 * 29 = 696
            10'b1100011110: z <= 10'b1011010000; // 24 * 30 = 720
            10'b1100011111: z <= 10'b1011101000; // 24 * 31 = 744
            10'b1100100000: z <= 10'b0000000000; // 25 * 0 = 0
            10'b1100100001: z <= 10'b0000011001; // 25 * 1 = 25
            10'b1100100010: z <= 10'b0000110010; // 25 * 2 = 50
            10'b1100100011: z <= 10'b0001001011; // 25 * 3 = 75
            10'b1100100100: z <= 10'b0001100100; // 25 * 4 = 100
            10'b1100100101: z <= 10'b0001111101; // 25 * 5 = 125
            10'b1100100110: z <= 10'b0010010110; // 25 * 6 = 150
            10'b1100100111: z <= 10'b0010101111; // 25 * 7 = 175
            10'b1100101000: z <= 10'b0011001000; // 25 * 8 = 200
            10'b1100101001: z <= 10'b0011100001; // 25 * 9 = 225
            10'b1100101010: z <= 10'b0011111010; // 25 * 10 = 250
            10'b1100101011: z <= 10'b0100010011; // 25 * 11 = 275
            10'b1100101100: z <= 10'b0100101100; // 25 * 12 = 300
            10'b1100101101: z <= 10'b0101000101; // 25 * 13 = 325
            10'b1100101110: z <= 10'b0101011110; // 25 * 14 = 350
            10'b1100101111: z <= 10'b0101110111; // 25 * 15 = 375
            10'b1100110000: z <= 10'b0110010000; // 25 * 16 = 400
            10'b1100110001: z <= 10'b0110101001; // 25 * 17 = 425
            10'b1100110010: z <= 10'b0111000010; // 25 * 18 = 450
            10'b1100110011: z <= 10'b0111011011; // 25 * 19 = 475
            10'b1100110100: z <= 10'b0111110100; // 25 * 20 = 500
            10'b1100110101: z <= 10'b1000001101; // 25 * 21 = 525
            10'b1100110110: z <= 10'b1000100110; // 25 * 22 = 550
            10'b1100110111: z <= 10'b1000111111; // 25 * 23 = 575
            10'b1100111000: z <= 10'b1001011000; // 25 * 24 = 600
            10'b1100111001: z <= 10'b1001110001; // 25 * 25 = 625
            10'b1100111010: z <= 10'b1010001010; // 25 * 26 = 650
            10'b1100111011: z <= 10'b1010100011; // 25 * 27 = 675
            10'b1100111100: z <= 10'b1010111100; // 25 * 28 = 700
            10'b1100111101: z <= 10'b1011010101; // 25 * 29 = 725
            10'b1100111110: z <= 10'b1011101110; // 25 * 30 = 750
            10'b1100111111: z <= 10'b1100000111; // 25 * 31 = 775
            10'b1101000000: z <= 10'b0000000000; // 26 * 0 = 0
            10'b1101000001: z <= 10'b0000011010; // 26 * 1 = 26
            10'b1101000010: z <= 10'b0000110100; // 26 * 2 = 52
            10'b1101000011: z <= 10'b0001001110; // 26 * 3 = 78
            10'b1101000100: z <= 10'b0001101000; // 26 * 4 = 104
            10'b1101000101: z <= 10'b0010000010; // 26 * 5 = 130
            10'b1101000110: z <= 10'b0010011100; // 26 * 6 = 156
            10'b1101000111: z <= 10'b0010110110; // 26 * 7 = 182
            10'b1101001000: z <= 10'b0011010000; // 26 * 8 = 208
            10'b1101001001: z <= 10'b0011101010; // 26 * 9 = 234
            10'b1101001010: z <= 10'b0100000100; // 26 * 10 = 260
            10'b1101001011: z <= 10'b0100011110; // 26 * 11 = 286
            10'b1101001100: z <= 10'b0100111000; // 26 * 12 = 312
            10'b1101001101: z <= 10'b0101010010; // 26 * 13 = 338
            10'b1101001110: z <= 10'b0101101100; // 26 * 14 = 364
            10'b1101001111: z <= 10'b0110000110; // 26 * 15 = 390
            10'b1101010000: z <= 10'b0110100000; // 26 * 16 = 416
            10'b1101010001: z <= 10'b0110111010; // 26 * 17 = 442
            10'b1101010010: z <= 10'b0111010100; // 26 * 18 = 468
            10'b1101010011: z <= 10'b0111101110; // 26 * 19 = 494
            10'b1101010100: z <= 10'b1000001000; // 26 * 20 = 520
            10'b1101010101: z <= 10'b1000100010; // 26 * 21 = 546
            10'b1101010110: z <= 10'b1000111100; // 26 * 22 = 572
            10'b1101010111: z <= 10'b1001010110; // 26 * 23 = 598
            10'b1101011000: z <= 10'b1001110000; // 26 * 24 = 624
            10'b1101011001: z <= 10'b1010001010; // 26 * 25 = 650
            10'b1101011010: z <= 10'b1010100100; // 26 * 26 = 676
            10'b1101011011: z <= 10'b1010111110; // 26 * 27 = 702
            10'b1101011100: z <= 10'b1011011000; // 26 * 28 = 728
            10'b1101011101: z <= 10'b1011110010; // 26 * 29 = 754
            10'b1101011110: z <= 10'b1100001100; // 26 * 30 = 780
            10'b1101011111: z <= 10'b1100100110; // 26 * 31 = 806
            10'b1101100000: z <= 10'b0000000000; // 27 * 0 = 0
            10'b1101100001: z <= 10'b0000011011; // 27 * 1 = 27
            10'b1101100010: z <= 10'b0000110110; // 27 * 2 = 54
            10'b1101100011: z <= 10'b0001010001; // 27 * 3 = 81
            10'b1101100100: z <= 10'b0001101100; // 27 * 4 = 108
            10'b1101100101: z <= 10'b0010000111; // 27 * 5 = 135
            10'b1101100110: z <= 10'b0010100010; // 27 * 6 = 162
            10'b1101100111: z <= 10'b0010111101; // 27 * 7 = 189
            10'b1101101000: z <= 10'b0011011000; // 27 * 8 = 216
            10'b1101101001: z <= 10'b0011110011; // 27 * 9 = 243
            10'b1101101010: z <= 10'b0100001110; // 27 * 10 = 270
            10'b1101101011: z <= 10'b0100101001; // 27 * 11 = 297
            10'b1101101100: z <= 10'b0101000100; // 27 * 12 = 324
            10'b1101101101: z <= 10'b0101011111; // 27 * 13 = 351
            10'b1101101110: z <= 10'b0101111010; // 27 * 14 = 378
            10'b1101101111: z <= 10'b0110010101; // 27 * 15 = 405
            10'b1101110000: z <= 10'b0110110000; // 27 * 16 = 432
            10'b1101110001: z <= 10'b0111001011; // 27 * 17 = 459
            10'b1101110010: z <= 10'b0111100110; // 27 * 18 = 486
            10'b1101110011: z <= 10'b1000000001; // 27 * 19 = 513
            10'b1101110100: z <= 10'b1000011100; // 27 * 20 = 540
            10'b1101110101: z <= 10'b1000110111; // 27 * 21 = 567
            10'b1101110110: z <= 10'b1001010010; // 27 * 22 = 594
            10'b1101110111: z <= 10'b1001101101; // 27 * 23 = 621
            10'b1101111000: z <= 10'b1010001000; // 27 * 24 = 648
            10'b1101111001: z <= 10'b1010100011; // 27 * 25 = 675
            10'b1101111010: z <= 10'b1010111110; // 27 * 26 = 702
            10'b1101111011: z <= 10'b1011011001; // 27 * 27 = 729
            10'b1101111100: z <= 10'b1011110100; // 27 * 28 = 756
            10'b1101111101: z <= 10'b1100001111; // 27 * 29 = 783
            10'b1101111110: z <= 10'b1100101010; // 27 * 30 = 810
            10'b1101111111: z <= 10'b1101000101; // 27 * 31 = 837
            10'b1110000000: z <= 10'b0000000000; // 28 * 0 = 0
            10'b1110000001: z <= 10'b0000011100; // 28 * 1 = 28
            10'b1110000010: z <= 10'b0000111000; // 28 * 2 = 56
            10'b1110000011: z <= 10'b0001010100; // 28 * 3 = 84
            10'b1110000100: z <= 10'b0001110000; // 28 * 4 = 112
            10'b1110000101: z <= 10'b0010001100; // 28 * 5 = 140
            10'b1110000110: z <= 10'b0010101000; // 28 * 6 = 168
            10'b1110000111: z <= 10'b0011000100; // 28 * 7 = 196
            10'b1110001000: z <= 10'b0011100000; // 28 * 8 = 224
            10'b1110001001: z <= 10'b0011111100; // 28 * 9 = 252
            10'b1110001010: z <= 10'b0100011000; // 28 * 10 = 280
            10'b1110001011: z <= 10'b0100110100; // 28 * 11 = 308
            10'b1110001100: z <= 10'b0101010000; // 28 * 12 = 336
            10'b1110001101: z <= 10'b0101101100; // 28 * 13 = 364
            10'b1110001110: z <= 10'b0110001000; // 28 * 14 = 392
            10'b1110001111: z <= 10'b0110100100; // 28 * 15 = 420
            10'b1110010000: z <= 10'b0111000000; // 28 * 16 = 448
            10'b1110010001: z <= 10'b0111011100; // 28 * 17 = 476
            10'b1110010010: z <= 10'b0111111000; // 28 * 18 = 504
            10'b1110010011: z <= 10'b1000010100; // 28 * 19 = 532
            10'b1110010100: z <= 10'b1000110000; // 28 * 20 = 560
            10'b1110010101: z <= 10'b1001001100; // 28 * 21 = 588
            10'b1110010110: z <= 10'b1001101000; // 28 * 22 = 616
            10'b1110010111: z <= 10'b1010000100; // 28 * 23 = 644
            10'b1110011000: z <= 10'b1010100000; // 28 * 24 = 672
            10'b1110011001: z <= 10'b1010111100; // 28 * 25 = 700
            10'b1110011010: z <= 10'b1011011000; // 28 * 26 = 728
            10'b1110011011: z <= 10'b1011110100; // 28 * 27 = 756
            10'b1110011100: z <= 10'b1100010000; // 28 * 28 = 784
            10'b1110011101: z <= 10'b1100101100; // 28 * 29 = 812
            10'b1110011110: z <= 10'b1101001000; // 28 * 30 = 840
            10'b1110011111: z <= 10'b1101100100; // 28 * 31 = 868
            10'b1110100000: z <= 10'b0000000000; // 29 * 0 = 0
            10'b1110100001: z <= 10'b0000011101; // 29 * 1 = 29
            10'b1110100010: z <= 10'b0000111010; // 29 * 2 = 58
            10'b1110100011: z <= 10'b0001010111; // 29 * 3 = 87
            10'b1110100100: z <= 10'b0001110100; // 29 * 4 = 116
            10'b1110100101: z <= 10'b0010010001; // 29 * 5 = 145
            10'b1110100110: z <= 10'b0010101110; // 29 * 6 = 174
            10'b1110100111: z <= 10'b0011001011; // 29 * 7 = 203
            10'b1110101000: z <= 10'b0011101000; // 29 * 8 = 232
            10'b1110101001: z <= 10'b0100000101; // 29 * 9 = 261
            10'b1110101010: z <= 10'b0100100010; // 29 * 10 = 290
            10'b1110101011: z <= 10'b0100111111; // 29 * 11 = 319
            10'b1110101100: z <= 10'b0101011100; // 29 * 12 = 348
            10'b1110101101: z <= 10'b0101111001; // 29 * 13 = 377
            10'b1110101110: z <= 10'b0110010110; // 29 * 14 = 406
            10'b1110101111: z <= 10'b0110110011; // 29 * 15 = 435
            10'b1110110000: z <= 10'b0111010000; // 29 * 16 = 464
            10'b1110110001: z <= 10'b0111101101; // 29 * 17 = 493
            10'b1110110010: z <= 10'b1000001010; // 29 * 18 = 522
            10'b1110110011: z <= 10'b1000100111; // 29 * 19 = 551
            10'b1110110100: z <= 10'b1001000100; // 29 * 20 = 580
            10'b1110110101: z <= 10'b1001100001; // 29 * 21 = 609
            10'b1110110110: z <= 10'b1001111110; // 29 * 22 = 638
            10'b1110110111: z <= 10'b1010011011; // 29 * 23 = 667
            10'b1110111000: z <= 10'b1010111000; // 29 * 24 = 696
            10'b1110111001: z <= 10'b1011010101; // 29 * 25 = 725
            10'b1110111010: z <= 10'b1011110010; // 29 * 26 = 754
            10'b1110111011: z <= 10'b1100001111; // 29 * 27 = 783
            10'b1110111100: z <= 10'b1100101100; // 29 * 28 = 812
            10'b1110111101: z <= 10'b1101001001; // 29 * 29 = 841
            10'b1110111110: z <= 10'b1101100110; // 29 * 30 = 870
            10'b1110111111: z <= 10'b1110000011; // 29 * 31 = 899
            10'b1111000000: z <= 10'b0000000000; // 30 * 0 = 0
            10'b1111000001: z <= 10'b0000011110; // 30 * 1 = 30
            10'b1111000010: z <= 10'b0000111100; // 30 * 2 = 60
            10'b1111000011: z <= 10'b0001011010; // 30 * 3 = 90
            10'b1111000100: z <= 10'b0001111000; // 30 * 4 = 120
            10'b1111000101: z <= 10'b0010010110; // 30 * 5 = 150
            10'b1111000110: z <= 10'b0010110100; // 30 * 6 = 180
            10'b1111000111: z <= 10'b0011010010; // 30 * 7 = 210
            10'b1111001000: z <= 10'b0011110000; // 30 * 8 = 240
            10'b1111001001: z <= 10'b0100001110; // 30 * 9 = 270
            10'b1111001010: z <= 10'b0100101100; // 30 * 10 = 300
            10'b1111001011: z <= 10'b0101001010; // 30 * 11 = 330
            10'b1111001100: z <= 10'b0101101000; // 30 * 12 = 360
            10'b1111001101: z <= 10'b0110000110; // 30 * 13 = 390
            10'b1111001110: z <= 10'b0110100100; // 30 * 14 = 420
            10'b1111001111: z <= 10'b0111000010; // 30 * 15 = 450
            10'b1111010000: z <= 10'b0111100000; // 30 * 16 = 480
            10'b1111010001: z <= 10'b0111111110; // 30 * 17 = 510
            10'b1111010010: z <= 10'b1000011100; // 30 * 18 = 540
            10'b1111010011: z <= 10'b1000111010; // 30 * 19 = 570
            10'b1111010100: z <= 10'b1001011000; // 30 * 20 = 600
            10'b1111010101: z <= 10'b1001110110; // 30 * 21 = 630
            10'b1111010110: z <= 10'b1010010100; // 30 * 22 = 660
            10'b1111010111: z <= 10'b1010110010; // 30 * 23 = 690
            10'b1111011000: z <= 10'b1011010000; // 30 * 24 = 720
            10'b1111011001: z <= 10'b1011101110; // 30 * 25 = 750
            10'b1111011010: z <= 10'b1100001100; // 30 * 26 = 780
            10'b1111011011: z <= 10'b1100101010; // 30 * 27 = 810
            10'b1111011100: z <= 10'b1101001000; // 30 * 28 = 840
            10'b1111011101: z <= 10'b1101100110; // 30 * 29 = 870
            10'b1111011110: z <= 10'b1110000100; // 30 * 30 = 900
            10'b1111011111: z <= 10'b1110100010; // 30 * 31 = 930
            10'b1111100000: z <= 10'b0000000000; // 31 * 0 = 0
            10'b1111100001: z <= 10'b0000011111; // 31 * 1 = 31
            10'b1111100010: z <= 10'b0000111110; // 31 * 2 = 62
            10'b1111100011: z <= 10'b0001011101; // 31 * 3 = 93
            10'b1111100100: z <= 10'b0001111100; // 31 * 4 = 124
            10'b1111100101: z <= 10'b0010011011; // 31 * 5 = 155
            10'b1111100110: z <= 10'b0010111010; // 31 * 6 = 186
            10'b1111100111: z <= 10'b0011011001; // 31 * 7 = 217
            10'b1111101000: z <= 10'b0011111000; // 31 * 8 = 248
            10'b1111101001: z <= 10'b0100010111; // 31 * 9 = 279
            10'b1111101010: z <= 10'b0100110110; // 31 * 10 = 310
            10'b1111101011: z <= 10'b0101010101; // 31 * 11 = 341
            10'b1111101100: z <= 10'b0101110100; // 31 * 12 = 372
            10'b1111101101: z <= 10'b0110010011; // 31 * 13 = 403
            10'b1111101110: z <= 10'b0110110010; // 31 * 14 = 434
            10'b1111101111: z <= 10'b0111010001; // 31 * 15 = 465
            10'b1111110000: z <= 10'b0111110000; // 31 * 16 = 496
            10'b1111110001: z <= 10'b1000001111; // 31 * 17 = 527
            10'b1111110010: z <= 10'b1000101110; // 31 * 18 = 558
            10'b1111110011: z <= 10'b1001001101; // 31 * 19 = 589
            10'b1111110100: z <= 10'b1001101100; // 31 * 20 = 620
            10'b1111110101: z <= 10'b1010001011; // 31 * 21 = 651
            10'b1111110110: z <= 10'b1010101010; // 31 * 22 = 682
            10'b1111110111: z <= 10'b1011001001; // 31 * 23 = 713
            10'b1111111000: z <= 10'b1011101000; // 31 * 24 = 744
            10'b1111111001: z <= 10'b1100000111; // 31 * 25 = 775
            10'b1111111010: z <= 10'b1100100110; // 31 * 26 = 806
            10'b1111111011: z <= 10'b1101000101; // 31 * 27 = 837
            10'b1111111100: z <= 10'b1101100100; // 31 * 28 = 868
            10'b1111111101: z <= 10'b1110000011; // 31 * 29 = 899
            10'b1111111110: z <= 10'b1110100010; // 31 * 30 = 930
            10'b1111111111: z <= 10'b1111000001; // 31 * 31 = 961
            default: z <= 0;
        endcase
        
    end


endmodule

